// http://www.ece.lsu.edu/ee3755/2002/l07.html

module s6bitdivider(q, r, a, b);
   input [5:0] a, b;

   output [5:0] q, r;

assign q[5] = 1'b0;
assign q[4] = ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0]));
assign q[3] = ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0]));
assign q[2] = ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0]));
assign q[1] = ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0]));
assign q[0] = ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0]));
assign r[5] = 1'b0;
assign r[4] = ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0]));
assign r[3] = ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0]));
assign r[2] = ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0]));
assign r[1] = ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0]));
assign r[0] = ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&(~a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&(~a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&(~a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&(~a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&(~a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&(~b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&(~b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&(~b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&(~b[4])&( b[3])&( b[2])&( b[1])&( b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&(~b[3])&( b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&(~b[2])&( b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&(~b[1])&(~b[0])) | ((~a[5])&( a[4])&( a[3])&( a[2])&( a[1])&( a[0])&(~b[5])&( b[4])&( b[3])&( b[2])&( b[1])&(~b[0]));
   endmodule
